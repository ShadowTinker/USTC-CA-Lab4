
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h28ce5d8c;
    ram_cell[       1] = 32'h0;  // 32'h705eac1b;
    ram_cell[       2] = 32'h0;  // 32'h61867afd;
    ram_cell[       3] = 32'h0;  // 32'ha9c7f5b0;
    ram_cell[       4] = 32'h0;  // 32'h02d2ecbb;
    ram_cell[       5] = 32'h0;  // 32'h2c748a56;
    ram_cell[       6] = 32'h0;  // 32'h09bc7e56;
    ram_cell[       7] = 32'h0;  // 32'h562676db;
    ram_cell[       8] = 32'h0;  // 32'h652ce53d;
    ram_cell[       9] = 32'h0;  // 32'h3a840d8f;
    ram_cell[      10] = 32'h0;  // 32'h014019aa;
    ram_cell[      11] = 32'h0;  // 32'h6f76fe3b;
    ram_cell[      12] = 32'h0;  // 32'h5826948a;
    ram_cell[      13] = 32'h0;  // 32'h75c1264e;
    ram_cell[      14] = 32'h0;  // 32'h20c2207a;
    ram_cell[      15] = 32'h0;  // 32'h84beea36;
    ram_cell[      16] = 32'h0;  // 32'h78f3cd78;
    ram_cell[      17] = 32'h0;  // 32'h7655de47;
    ram_cell[      18] = 32'h0;  // 32'h32ebd90e;
    ram_cell[      19] = 32'h0;  // 32'h0a81c255;
    ram_cell[      20] = 32'h0;  // 32'hf5b13f15;
    ram_cell[      21] = 32'h0;  // 32'hb01e4d1f;
    ram_cell[      22] = 32'h0;  // 32'h27cbd7fc;
    ram_cell[      23] = 32'h0;  // 32'h860f282b;
    ram_cell[      24] = 32'h0;  // 32'h1fcf4cfd;
    ram_cell[      25] = 32'h0;  // 32'hbf816ee8;
    ram_cell[      26] = 32'h0;  // 32'h2b50684e;
    ram_cell[      27] = 32'h0;  // 32'h438607e6;
    ram_cell[      28] = 32'h0;  // 32'hd7a7f4c9;
    ram_cell[      29] = 32'h0;  // 32'hdd4b7109;
    ram_cell[      30] = 32'h0;  // 32'h6e79c348;
    ram_cell[      31] = 32'h0;  // 32'hee2fb741;
    ram_cell[      32] = 32'h0;  // 32'hc2fde9bd;
    ram_cell[      33] = 32'h0;  // 32'ha3920453;
    ram_cell[      34] = 32'h0;  // 32'h4411789f;
    ram_cell[      35] = 32'h0;  // 32'h90216d80;
    ram_cell[      36] = 32'h0;  // 32'hb13f35fa;
    ram_cell[      37] = 32'h0;  // 32'hbf8edf00;
    ram_cell[      38] = 32'h0;  // 32'hf9c82204;
    ram_cell[      39] = 32'h0;  // 32'he15077f6;
    ram_cell[      40] = 32'h0;  // 32'had0144e0;
    ram_cell[      41] = 32'h0;  // 32'h4f14be22;
    ram_cell[      42] = 32'h0;  // 32'hcc749af2;
    ram_cell[      43] = 32'h0;  // 32'h104db8a2;
    ram_cell[      44] = 32'h0;  // 32'h66b6bd26;
    ram_cell[      45] = 32'h0;  // 32'he1452f33;
    ram_cell[      46] = 32'h0;  // 32'hcef536b6;
    ram_cell[      47] = 32'h0;  // 32'h1bfc1fbf;
    ram_cell[      48] = 32'h0;  // 32'h0b904559;
    ram_cell[      49] = 32'h0;  // 32'hffbbb18f;
    ram_cell[      50] = 32'h0;  // 32'hff77f1ef;
    ram_cell[      51] = 32'h0;  // 32'hb2984412;
    ram_cell[      52] = 32'h0;  // 32'hba281738;
    ram_cell[      53] = 32'h0;  // 32'he4c074a4;
    ram_cell[      54] = 32'h0;  // 32'hebf3bddf;
    ram_cell[      55] = 32'h0;  // 32'hbc25efdf;
    ram_cell[      56] = 32'h0;  // 32'h959a03ee;
    ram_cell[      57] = 32'h0;  // 32'h88b7d444;
    ram_cell[      58] = 32'h0;  // 32'h918f692c;
    ram_cell[      59] = 32'h0;  // 32'h15ad1851;
    ram_cell[      60] = 32'h0;  // 32'h354e0bbd;
    ram_cell[      61] = 32'h0;  // 32'hdff87d94;
    ram_cell[      62] = 32'h0;  // 32'h08410a3d;
    ram_cell[      63] = 32'h0;  // 32'hdf19b8d7;
    ram_cell[      64] = 32'h0;  // 32'h29bf647e;
    ram_cell[      65] = 32'h0;  // 32'hca7d30a3;
    ram_cell[      66] = 32'h0;  // 32'hde54c411;
    ram_cell[      67] = 32'h0;  // 32'hf33f92df;
    ram_cell[      68] = 32'h0;  // 32'had088ce6;
    ram_cell[      69] = 32'h0;  // 32'h08d9fe1f;
    ram_cell[      70] = 32'h0;  // 32'hb6aae3ce;
    ram_cell[      71] = 32'h0;  // 32'hfd202896;
    ram_cell[      72] = 32'h0;  // 32'h5e2ac290;
    ram_cell[      73] = 32'h0;  // 32'he6110509;
    ram_cell[      74] = 32'h0;  // 32'h97eab454;
    ram_cell[      75] = 32'h0;  // 32'hbdb0b46d;
    ram_cell[      76] = 32'h0;  // 32'he4f9dcde;
    ram_cell[      77] = 32'h0;  // 32'h28fabf24;
    ram_cell[      78] = 32'h0;  // 32'h72a8d46c;
    ram_cell[      79] = 32'h0;  // 32'h6aa77543;
    ram_cell[      80] = 32'h0;  // 32'h41bd1d2b;
    ram_cell[      81] = 32'h0;  // 32'h0e03bb6c;
    ram_cell[      82] = 32'h0;  // 32'hcb951970;
    ram_cell[      83] = 32'h0;  // 32'h41a411c5;
    ram_cell[      84] = 32'h0;  // 32'h180f9a96;
    ram_cell[      85] = 32'h0;  // 32'hba285bc1;
    ram_cell[      86] = 32'h0;  // 32'h5c13e266;
    ram_cell[      87] = 32'h0;  // 32'h37224660;
    ram_cell[      88] = 32'h0;  // 32'h22984b8b;
    ram_cell[      89] = 32'h0;  // 32'h7e665c2d;
    ram_cell[      90] = 32'h0;  // 32'h77706dd9;
    ram_cell[      91] = 32'h0;  // 32'h38f6d3c7;
    ram_cell[      92] = 32'h0;  // 32'h56556847;
    ram_cell[      93] = 32'h0;  // 32'hcad20745;
    ram_cell[      94] = 32'h0;  // 32'h30827524;
    ram_cell[      95] = 32'h0;  // 32'ha3088694;
    ram_cell[      96] = 32'h0;  // 32'h4072838a;
    ram_cell[      97] = 32'h0;  // 32'hf1f3f2d7;
    ram_cell[      98] = 32'h0;  // 32'h8cc6585f;
    ram_cell[      99] = 32'h0;  // 32'hcf893e3f;
    ram_cell[     100] = 32'h0;  // 32'h84f06f25;
    ram_cell[     101] = 32'h0;  // 32'h91baff73;
    ram_cell[     102] = 32'h0;  // 32'h64a6694f;
    ram_cell[     103] = 32'h0;  // 32'hcbfebab5;
    ram_cell[     104] = 32'h0;  // 32'hc2f55aa3;
    ram_cell[     105] = 32'h0;  // 32'h4454c7e2;
    ram_cell[     106] = 32'h0;  // 32'h452bdfc9;
    ram_cell[     107] = 32'h0;  // 32'h9591e698;
    ram_cell[     108] = 32'h0;  // 32'h2088ccb7;
    ram_cell[     109] = 32'h0;  // 32'h49e74ed3;
    ram_cell[     110] = 32'h0;  // 32'hbce2e34f;
    ram_cell[     111] = 32'h0;  // 32'hac860a3d;
    ram_cell[     112] = 32'h0;  // 32'h0e475299;
    ram_cell[     113] = 32'h0;  // 32'h8130bac8;
    ram_cell[     114] = 32'h0;  // 32'hc51c5a98;
    ram_cell[     115] = 32'h0;  // 32'h6e565900;
    ram_cell[     116] = 32'h0;  // 32'h7435e4eb;
    ram_cell[     117] = 32'h0;  // 32'ha3825edf;
    ram_cell[     118] = 32'h0;  // 32'hbf176dfa;
    ram_cell[     119] = 32'h0;  // 32'hd047d5a3;
    ram_cell[     120] = 32'h0;  // 32'h25374905;
    ram_cell[     121] = 32'h0;  // 32'hd5220298;
    ram_cell[     122] = 32'h0;  // 32'hffbc5365;
    ram_cell[     123] = 32'h0;  // 32'h1f8cf632;
    ram_cell[     124] = 32'h0;  // 32'hbc410ad6;
    ram_cell[     125] = 32'h0;  // 32'he3a2779e;
    ram_cell[     126] = 32'h0;  // 32'h642e9aa3;
    ram_cell[     127] = 32'h0;  // 32'hd430832d;
    ram_cell[     128] = 32'h0;  // 32'h000a12e9;
    ram_cell[     129] = 32'h0;  // 32'h6c7dc2e9;
    ram_cell[     130] = 32'h0;  // 32'h85210671;
    ram_cell[     131] = 32'h0;  // 32'h3a0e760f;
    ram_cell[     132] = 32'h0;  // 32'h0bef0d2d;
    ram_cell[     133] = 32'h0;  // 32'h392a4e9f;
    ram_cell[     134] = 32'h0;  // 32'hd8b982a5;
    ram_cell[     135] = 32'h0;  // 32'h45eb4342;
    ram_cell[     136] = 32'h0;  // 32'h0064305b;
    ram_cell[     137] = 32'h0;  // 32'h942eebc6;
    ram_cell[     138] = 32'h0;  // 32'ha6d7cf8f;
    ram_cell[     139] = 32'h0;  // 32'h688c8a09;
    ram_cell[     140] = 32'h0;  // 32'h08375a49;
    ram_cell[     141] = 32'h0;  // 32'hcd7efaca;
    ram_cell[     142] = 32'h0;  // 32'haddedef9;
    ram_cell[     143] = 32'h0;  // 32'he485a0c7;
    ram_cell[     144] = 32'h0;  // 32'hd95ba9a6;
    ram_cell[     145] = 32'h0;  // 32'hfac42bc0;
    ram_cell[     146] = 32'h0;  // 32'h1a9410ab;
    ram_cell[     147] = 32'h0;  // 32'h90373f37;
    ram_cell[     148] = 32'h0;  // 32'h672e0389;
    ram_cell[     149] = 32'h0;  // 32'hca79476e;
    ram_cell[     150] = 32'h0;  // 32'h6c1b583a;
    ram_cell[     151] = 32'h0;  // 32'hd3a75d6e;
    ram_cell[     152] = 32'h0;  // 32'h83382911;
    ram_cell[     153] = 32'h0;  // 32'h53e1d323;
    ram_cell[     154] = 32'h0;  // 32'h2faf03c3;
    ram_cell[     155] = 32'h0;  // 32'h21fc3b36;
    ram_cell[     156] = 32'h0;  // 32'h57b374f7;
    ram_cell[     157] = 32'h0;  // 32'h67105662;
    ram_cell[     158] = 32'h0;  // 32'h17e66c34;
    ram_cell[     159] = 32'h0;  // 32'hb2cc1467;
    ram_cell[     160] = 32'h0;  // 32'h72fb6646;
    ram_cell[     161] = 32'h0;  // 32'hf8006670;
    ram_cell[     162] = 32'h0;  // 32'h84455c8e;
    ram_cell[     163] = 32'h0;  // 32'h9d6ed0da;
    ram_cell[     164] = 32'h0;  // 32'hecc97d67;
    ram_cell[     165] = 32'h0;  // 32'hdb2ec7bc;
    ram_cell[     166] = 32'h0;  // 32'h539a5aaa;
    ram_cell[     167] = 32'h0;  // 32'h54dfeaf7;
    ram_cell[     168] = 32'h0;  // 32'hf1128b77;
    ram_cell[     169] = 32'h0;  // 32'hab51d3e8;
    ram_cell[     170] = 32'h0;  // 32'hbe5fcbf2;
    ram_cell[     171] = 32'h0;  // 32'h1b4582f9;
    ram_cell[     172] = 32'h0;  // 32'h560ca596;
    ram_cell[     173] = 32'h0;  // 32'h5e98fe54;
    ram_cell[     174] = 32'h0;  // 32'h7d9c2e55;
    ram_cell[     175] = 32'h0;  // 32'h91f0e63c;
    ram_cell[     176] = 32'h0;  // 32'h4bb96d97;
    ram_cell[     177] = 32'h0;  // 32'hcbe33a22;
    ram_cell[     178] = 32'h0;  // 32'h521840d5;
    ram_cell[     179] = 32'h0;  // 32'h49861126;
    ram_cell[     180] = 32'h0;  // 32'h19b34a36;
    ram_cell[     181] = 32'h0;  // 32'h365d1bfb;
    ram_cell[     182] = 32'h0;  // 32'hc12e1ed7;
    ram_cell[     183] = 32'h0;  // 32'h24a4c44b;
    ram_cell[     184] = 32'h0;  // 32'hf9b51386;
    ram_cell[     185] = 32'h0;  // 32'h35ae43aa;
    ram_cell[     186] = 32'h0;  // 32'hac5b1b56;
    ram_cell[     187] = 32'h0;  // 32'h26d7f379;
    ram_cell[     188] = 32'h0;  // 32'h49f78925;
    ram_cell[     189] = 32'h0;  // 32'hdb052fa2;
    ram_cell[     190] = 32'h0;  // 32'h461d003e;
    ram_cell[     191] = 32'h0;  // 32'hd10c81c5;
    ram_cell[     192] = 32'h0;  // 32'h0f747b25;
    ram_cell[     193] = 32'h0;  // 32'h60f4bed6;
    ram_cell[     194] = 32'h0;  // 32'h42ec3682;
    ram_cell[     195] = 32'h0;  // 32'h33df3e18;
    ram_cell[     196] = 32'h0;  // 32'hfd343ae4;
    ram_cell[     197] = 32'h0;  // 32'h3b94f8b1;
    ram_cell[     198] = 32'h0;  // 32'h7fc54a3b;
    ram_cell[     199] = 32'h0;  // 32'h0c009d73;
    ram_cell[     200] = 32'h0;  // 32'hfc54295a;
    ram_cell[     201] = 32'h0;  // 32'hab3b9a69;
    ram_cell[     202] = 32'h0;  // 32'hab3697fe;
    ram_cell[     203] = 32'h0;  // 32'hb14c27c3;
    ram_cell[     204] = 32'h0;  // 32'h829fda82;
    ram_cell[     205] = 32'h0;  // 32'had394a28;
    ram_cell[     206] = 32'h0;  // 32'h776cae13;
    ram_cell[     207] = 32'h0;  // 32'hb0476999;
    ram_cell[     208] = 32'h0;  // 32'h603f1c45;
    ram_cell[     209] = 32'h0;  // 32'hf47d5d7d;
    ram_cell[     210] = 32'h0;  // 32'h417d0fb1;
    ram_cell[     211] = 32'h0;  // 32'h006b33d1;
    ram_cell[     212] = 32'h0;  // 32'h173ca34d;
    ram_cell[     213] = 32'h0;  // 32'h96b8e4fb;
    ram_cell[     214] = 32'h0;  // 32'hb20211b2;
    ram_cell[     215] = 32'h0;  // 32'hd6159d90;
    ram_cell[     216] = 32'h0;  // 32'h8c53cd06;
    ram_cell[     217] = 32'h0;  // 32'hdb0c72b1;
    ram_cell[     218] = 32'h0;  // 32'h106e9e03;
    ram_cell[     219] = 32'h0;  // 32'h6f883f04;
    ram_cell[     220] = 32'h0;  // 32'h02e0b5ff;
    ram_cell[     221] = 32'h0;  // 32'hd94c9f79;
    ram_cell[     222] = 32'h0;  // 32'hef55c8a7;
    ram_cell[     223] = 32'h0;  // 32'hc0efb598;
    ram_cell[     224] = 32'h0;  // 32'h09471463;
    ram_cell[     225] = 32'h0;  // 32'h588a8cf0;
    ram_cell[     226] = 32'h0;  // 32'h9cb2ed11;
    ram_cell[     227] = 32'h0;  // 32'hff58a9f4;
    ram_cell[     228] = 32'h0;  // 32'h44adcab1;
    ram_cell[     229] = 32'h0;  // 32'h47ac4fa0;
    ram_cell[     230] = 32'h0;  // 32'h20f5987e;
    ram_cell[     231] = 32'h0;  // 32'h4c152446;
    ram_cell[     232] = 32'h0;  // 32'h612dc2f1;
    ram_cell[     233] = 32'h0;  // 32'he491fa24;
    ram_cell[     234] = 32'h0;  // 32'hd9286bc5;
    ram_cell[     235] = 32'h0;  // 32'h98905876;
    ram_cell[     236] = 32'h0;  // 32'hefefeb0e;
    ram_cell[     237] = 32'h0;  // 32'h69703eaf;
    ram_cell[     238] = 32'h0;  // 32'hd97b3c58;
    ram_cell[     239] = 32'h0;  // 32'h0f9a777b;
    ram_cell[     240] = 32'h0;  // 32'ha11819a6;
    ram_cell[     241] = 32'h0;  // 32'h6e1c6541;
    ram_cell[     242] = 32'h0;  // 32'h54430668;
    ram_cell[     243] = 32'h0;  // 32'h1e096979;
    ram_cell[     244] = 32'h0;  // 32'hbc101f8d;
    ram_cell[     245] = 32'h0;  // 32'hec611371;
    ram_cell[     246] = 32'h0;  // 32'h7efb2e39;
    ram_cell[     247] = 32'h0;  // 32'ha7bb438a;
    ram_cell[     248] = 32'h0;  // 32'h36fc2cc5;
    ram_cell[     249] = 32'h0;  // 32'hd3455746;
    ram_cell[     250] = 32'h0;  // 32'h345d9db0;
    ram_cell[     251] = 32'h0;  // 32'h5320fa36;
    ram_cell[     252] = 32'h0;  // 32'hfc2501b0;
    ram_cell[     253] = 32'h0;  // 32'h268a61eb;
    ram_cell[     254] = 32'h0;  // 32'hd5ea83e6;
    ram_cell[     255] = 32'h0;  // 32'h93209397;
    // src matrix A
    ram_cell[     256] = 32'h02fef0ab;
    ram_cell[     257] = 32'h50ca985f;
    ram_cell[     258] = 32'h1069bc69;
    ram_cell[     259] = 32'hed19e344;
    ram_cell[     260] = 32'h3bd85ef2;
    ram_cell[     261] = 32'hc3ce5b7a;
    ram_cell[     262] = 32'hc383b1c1;
    ram_cell[     263] = 32'h5555a29a;
    ram_cell[     264] = 32'h086534f8;
    ram_cell[     265] = 32'h0f47c348;
    ram_cell[     266] = 32'h9137decc;
    ram_cell[     267] = 32'h682a10bc;
    ram_cell[     268] = 32'h9ace8fdd;
    ram_cell[     269] = 32'he65ce047;
    ram_cell[     270] = 32'h0c620550;
    ram_cell[     271] = 32'he993a1c0;
    ram_cell[     272] = 32'h9d258088;
    ram_cell[     273] = 32'h61088748;
    ram_cell[     274] = 32'hdf652ce2;
    ram_cell[     275] = 32'h87f26ff5;
    ram_cell[     276] = 32'h39cfb031;
    ram_cell[     277] = 32'hce648b5b;
    ram_cell[     278] = 32'he95017b1;
    ram_cell[     279] = 32'hbc319ec5;
    ram_cell[     280] = 32'h4fe10e3c;
    ram_cell[     281] = 32'ha599e327;
    ram_cell[     282] = 32'he2d9849c;
    ram_cell[     283] = 32'h7cf11a50;
    ram_cell[     284] = 32'h47ff0777;
    ram_cell[     285] = 32'h6e552e42;
    ram_cell[     286] = 32'hfe2804de;
    ram_cell[     287] = 32'h648bd393;
    ram_cell[     288] = 32'h756f9cec;
    ram_cell[     289] = 32'hfc2d96ef;
    ram_cell[     290] = 32'ha02afc30;
    ram_cell[     291] = 32'h1ade0255;
    ram_cell[     292] = 32'h77bfdbdb;
    ram_cell[     293] = 32'hd872ca3f;
    ram_cell[     294] = 32'h9e5213b2;
    ram_cell[     295] = 32'hc5407072;
    ram_cell[     296] = 32'hd6ad1815;
    ram_cell[     297] = 32'h59f9c589;
    ram_cell[     298] = 32'h10c4ccbf;
    ram_cell[     299] = 32'h1d4bec86;
    ram_cell[     300] = 32'ha6e25b92;
    ram_cell[     301] = 32'he7db1227;
    ram_cell[     302] = 32'h3d00cb52;
    ram_cell[     303] = 32'h1f98bc28;
    ram_cell[     304] = 32'hdb9ca56d;
    ram_cell[     305] = 32'h4c4c555d;
    ram_cell[     306] = 32'hd74698e1;
    ram_cell[     307] = 32'haa5dadfd;
    ram_cell[     308] = 32'hbc5b9fd0;
    ram_cell[     309] = 32'h7c742397;
    ram_cell[     310] = 32'hbd038e6c;
    ram_cell[     311] = 32'he38208f8;
    ram_cell[     312] = 32'hd9ae91a1;
    ram_cell[     313] = 32'h0e1d2129;
    ram_cell[     314] = 32'hc7722223;
    ram_cell[     315] = 32'ha5c56cce;
    ram_cell[     316] = 32'hf8c8a4ec;
    ram_cell[     317] = 32'h74e3395a;
    ram_cell[     318] = 32'h85689fc2;
    ram_cell[     319] = 32'h050d5b7f;
    ram_cell[     320] = 32'h5acffdcf;
    ram_cell[     321] = 32'h44badd21;
    ram_cell[     322] = 32'h6743bae5;
    ram_cell[     323] = 32'hc08b6f1c;
    ram_cell[     324] = 32'h873d4d2c;
    ram_cell[     325] = 32'hfda081d6;
    ram_cell[     326] = 32'h3e8bf065;
    ram_cell[     327] = 32'he1e068c6;
    ram_cell[     328] = 32'h596507b9;
    ram_cell[     329] = 32'h6de399b9;
    ram_cell[     330] = 32'h1cfc4989;
    ram_cell[     331] = 32'h1bbba6b0;
    ram_cell[     332] = 32'ha7682287;
    ram_cell[     333] = 32'h40c48692;
    ram_cell[     334] = 32'h0df1a55c;
    ram_cell[     335] = 32'hf7cdae45;
    ram_cell[     336] = 32'he45658f1;
    ram_cell[     337] = 32'h4d72fc14;
    ram_cell[     338] = 32'hc3126102;
    ram_cell[     339] = 32'h33f0d5d3;
    ram_cell[     340] = 32'he7d125ee;
    ram_cell[     341] = 32'hc1602a2a;
    ram_cell[     342] = 32'h8bd289b1;
    ram_cell[     343] = 32'h783c1520;
    ram_cell[     344] = 32'h2229f4ad;
    ram_cell[     345] = 32'hc416f831;
    ram_cell[     346] = 32'h7f066b2a;
    ram_cell[     347] = 32'h516e04f1;
    ram_cell[     348] = 32'hd647050a;
    ram_cell[     349] = 32'hbe6958d3;
    ram_cell[     350] = 32'hffff02d9;
    ram_cell[     351] = 32'hd6c4d81c;
    ram_cell[     352] = 32'h28966581;
    ram_cell[     353] = 32'h690353cf;
    ram_cell[     354] = 32'h709cb66e;
    ram_cell[     355] = 32'h31a893c2;
    ram_cell[     356] = 32'ha732a3c9;
    ram_cell[     357] = 32'h12593985;
    ram_cell[     358] = 32'h2f679c0e;
    ram_cell[     359] = 32'he7c489a6;
    ram_cell[     360] = 32'h90d671bf;
    ram_cell[     361] = 32'hbd50e2f9;
    ram_cell[     362] = 32'hd7d1c4dc;
    ram_cell[     363] = 32'h1bea76f8;
    ram_cell[     364] = 32'h06fba261;
    ram_cell[     365] = 32'hdecfe4eb;
    ram_cell[     366] = 32'h02addeca;
    ram_cell[     367] = 32'ha1c9a781;
    ram_cell[     368] = 32'hae421364;
    ram_cell[     369] = 32'hedeba803;
    ram_cell[     370] = 32'h0e5011d6;
    ram_cell[     371] = 32'hb66058e2;
    ram_cell[     372] = 32'h9055f00b;
    ram_cell[     373] = 32'h74de2ca1;
    ram_cell[     374] = 32'h72dd4b07;
    ram_cell[     375] = 32'h58066055;
    ram_cell[     376] = 32'h74140d4f;
    ram_cell[     377] = 32'hd651a914;
    ram_cell[     378] = 32'h2315331f;
    ram_cell[     379] = 32'h49e84d91;
    ram_cell[     380] = 32'h7c835142;
    ram_cell[     381] = 32'hffe411fd;
    ram_cell[     382] = 32'h7fd8e84a;
    ram_cell[     383] = 32'ha2e5f87a;
    ram_cell[     384] = 32'hfa6cbf65;
    ram_cell[     385] = 32'h2aed1b05;
    ram_cell[     386] = 32'h7ca3563e;
    ram_cell[     387] = 32'h42b20d59;
    ram_cell[     388] = 32'h91fb6d19;
    ram_cell[     389] = 32'h315f37a4;
    ram_cell[     390] = 32'hb92e0779;
    ram_cell[     391] = 32'h5145508f;
    ram_cell[     392] = 32'h5db4ccd9;
    ram_cell[     393] = 32'hb1eacd07;
    ram_cell[     394] = 32'hbc034e30;
    ram_cell[     395] = 32'hcab4c133;
    ram_cell[     396] = 32'h84591661;
    ram_cell[     397] = 32'h0a94bb70;
    ram_cell[     398] = 32'h0e1f3811;
    ram_cell[     399] = 32'h028fd49b;
    ram_cell[     400] = 32'h31e7c509;
    ram_cell[     401] = 32'he1acf370;
    ram_cell[     402] = 32'h2b5fa277;
    ram_cell[     403] = 32'h299496f8;
    ram_cell[     404] = 32'h3674b4bf;
    ram_cell[     405] = 32'h61234415;
    ram_cell[     406] = 32'hd2133d7f;
    ram_cell[     407] = 32'h2bd1d78d;
    ram_cell[     408] = 32'h5984f2d4;
    ram_cell[     409] = 32'h4a525379;
    ram_cell[     410] = 32'hd855ed70;
    ram_cell[     411] = 32'h4925bcb6;
    ram_cell[     412] = 32'hdf5986b6;
    ram_cell[     413] = 32'h935ccf20;
    ram_cell[     414] = 32'h1cc0b315;
    ram_cell[     415] = 32'h2727ed27;
    ram_cell[     416] = 32'h310991c6;
    ram_cell[     417] = 32'h1c99cb80;
    ram_cell[     418] = 32'ha8bd5d57;
    ram_cell[     419] = 32'h08f17293;
    ram_cell[     420] = 32'hd3e0a1fc;
    ram_cell[     421] = 32'h41f385ea;
    ram_cell[     422] = 32'h90b24936;
    ram_cell[     423] = 32'h56555abc;
    ram_cell[     424] = 32'h9349e000;
    ram_cell[     425] = 32'h5c91b436;
    ram_cell[     426] = 32'hffadd078;
    ram_cell[     427] = 32'hbca394a6;
    ram_cell[     428] = 32'h4d7bf8a7;
    ram_cell[     429] = 32'h38e68767;
    ram_cell[     430] = 32'he27d7434;
    ram_cell[     431] = 32'ha2c8d16b;
    ram_cell[     432] = 32'hec45430a;
    ram_cell[     433] = 32'h1c1194ee;
    ram_cell[     434] = 32'h9d03b742;
    ram_cell[     435] = 32'he195ecdb;
    ram_cell[     436] = 32'h35c9c4e9;
    ram_cell[     437] = 32'h62271340;
    ram_cell[     438] = 32'h4d01a91a;
    ram_cell[     439] = 32'h4ed2b103;
    ram_cell[     440] = 32'h8b0830c5;
    ram_cell[     441] = 32'h0847567f;
    ram_cell[     442] = 32'ha963579c;
    ram_cell[     443] = 32'h0bcfe8d5;
    ram_cell[     444] = 32'h2f3010c6;
    ram_cell[     445] = 32'hb270ed1c;
    ram_cell[     446] = 32'h14c5db43;
    ram_cell[     447] = 32'h44bc5cfe;
    ram_cell[     448] = 32'h09b60a96;
    ram_cell[     449] = 32'had179c21;
    ram_cell[     450] = 32'ha6ccc742;
    ram_cell[     451] = 32'h9c45614d;
    ram_cell[     452] = 32'h747a2d95;
    ram_cell[     453] = 32'h56514bd9;
    ram_cell[     454] = 32'h4de33bd9;
    ram_cell[     455] = 32'h255e33d0;
    ram_cell[     456] = 32'ha9b85565;
    ram_cell[     457] = 32'h917c2a3b;
    ram_cell[     458] = 32'h10b0f06b;
    ram_cell[     459] = 32'h6d4c19f8;
    ram_cell[     460] = 32'h30d6e695;
    ram_cell[     461] = 32'hf7aa41f3;
    ram_cell[     462] = 32'h8e76d81c;
    ram_cell[     463] = 32'hda334a87;
    ram_cell[     464] = 32'hf5829b86;
    ram_cell[     465] = 32'h0a969a11;
    ram_cell[     466] = 32'h2081776a;
    ram_cell[     467] = 32'h35adb857;
    ram_cell[     468] = 32'h593d28fe;
    ram_cell[     469] = 32'he681eeae;
    ram_cell[     470] = 32'h50e91d78;
    ram_cell[     471] = 32'h2c799812;
    ram_cell[     472] = 32'h437b0105;
    ram_cell[     473] = 32'hd31576a6;
    ram_cell[     474] = 32'h3d2c0f3d;
    ram_cell[     475] = 32'h86576c64;
    ram_cell[     476] = 32'hac4a8103;
    ram_cell[     477] = 32'h0f34e0bb;
    ram_cell[     478] = 32'h3467704b;
    ram_cell[     479] = 32'h4109abe2;
    ram_cell[     480] = 32'h656ac54f;
    ram_cell[     481] = 32'h091cea2f;
    ram_cell[     482] = 32'h99adc8a8;
    ram_cell[     483] = 32'h6995c999;
    ram_cell[     484] = 32'hc2a8e6d1;
    ram_cell[     485] = 32'h2ba47e44;
    ram_cell[     486] = 32'hb76b9fe9;
    ram_cell[     487] = 32'h67c02c90;
    ram_cell[     488] = 32'hd4ff2312;
    ram_cell[     489] = 32'h1ee49d3f;
    ram_cell[     490] = 32'h6a36771b;
    ram_cell[     491] = 32'hf6d9af16;
    ram_cell[     492] = 32'hf83268f4;
    ram_cell[     493] = 32'h353b32fa;
    ram_cell[     494] = 32'h557ab592;
    ram_cell[     495] = 32'h4e7cc164;
    ram_cell[     496] = 32'h91706453;
    ram_cell[     497] = 32'h43d4d275;
    ram_cell[     498] = 32'hb5169d1f;
    ram_cell[     499] = 32'ha4f73025;
    ram_cell[     500] = 32'h319877d3;
    ram_cell[     501] = 32'h0b3c8cdd;
    ram_cell[     502] = 32'hbfc49f64;
    ram_cell[     503] = 32'h12a71dcb;
    ram_cell[     504] = 32'hd1fa8b16;
    ram_cell[     505] = 32'hd416ca93;
    ram_cell[     506] = 32'h8fcb5f25;
    ram_cell[     507] = 32'h3c062c6d;
    ram_cell[     508] = 32'h75a59da6;
    ram_cell[     509] = 32'h004a2eaf;
    ram_cell[     510] = 32'h56cf8627;
    ram_cell[     511] = 32'hef08444b;
    // src matrix B
    ram_cell[     512] = 32'ha76463fd;
    ram_cell[     513] = 32'he7066734;
    ram_cell[     514] = 32'hafe72327;
    ram_cell[     515] = 32'hd68dfd2d;
    ram_cell[     516] = 32'ha05bd0bd;
    ram_cell[     517] = 32'hcce559eb;
    ram_cell[     518] = 32'h9e03e36e;
    ram_cell[     519] = 32'hd3c7da71;
    ram_cell[     520] = 32'h90ec65d6;
    ram_cell[     521] = 32'h21a676cc;
    ram_cell[     522] = 32'h4da7ee5e;
    ram_cell[     523] = 32'hb107d9e7;
    ram_cell[     524] = 32'h878472f0;
    ram_cell[     525] = 32'hb1ee8958;
    ram_cell[     526] = 32'h0b190ce3;
    ram_cell[     527] = 32'h0b853697;
    ram_cell[     528] = 32'h924c4ef9;
    ram_cell[     529] = 32'h750ade3a;
    ram_cell[     530] = 32'h4d296f1a;
    ram_cell[     531] = 32'h16872414;
    ram_cell[     532] = 32'h0bb64ec4;
    ram_cell[     533] = 32'h2b2ca5a2;
    ram_cell[     534] = 32'hfd211291;
    ram_cell[     535] = 32'h9388b0cb;
    ram_cell[     536] = 32'h8486ae61;
    ram_cell[     537] = 32'h50a618ad;
    ram_cell[     538] = 32'hd6a51f4d;
    ram_cell[     539] = 32'hfbcbc36e;
    ram_cell[     540] = 32'h5fef967a;
    ram_cell[     541] = 32'h159819fd;
    ram_cell[     542] = 32'ha14ae1f3;
    ram_cell[     543] = 32'hb78cf629;
    ram_cell[     544] = 32'h1fc749fc;
    ram_cell[     545] = 32'hc0e540da;
    ram_cell[     546] = 32'ha4bb3710;
    ram_cell[     547] = 32'h90b0bb77;
    ram_cell[     548] = 32'h8509f900;
    ram_cell[     549] = 32'h75e41a07;
    ram_cell[     550] = 32'h56defa8a;
    ram_cell[     551] = 32'h7abfc884;
    ram_cell[     552] = 32'ha6dec095;
    ram_cell[     553] = 32'h3b818ab7;
    ram_cell[     554] = 32'hcac64389;
    ram_cell[     555] = 32'heee57aca;
    ram_cell[     556] = 32'h4253ab5d;
    ram_cell[     557] = 32'h446bac43;
    ram_cell[     558] = 32'h7d8094f9;
    ram_cell[     559] = 32'h5c18f6b2;
    ram_cell[     560] = 32'h1469960b;
    ram_cell[     561] = 32'h6c34c6ca;
    ram_cell[     562] = 32'h3dc08e16;
    ram_cell[     563] = 32'h9b97e81f;
    ram_cell[     564] = 32'ha30d6696;
    ram_cell[     565] = 32'hb669fad4;
    ram_cell[     566] = 32'hf54b316e;
    ram_cell[     567] = 32'hc4995f4c;
    ram_cell[     568] = 32'h8a5503ff;
    ram_cell[     569] = 32'h5989142c;
    ram_cell[     570] = 32'h12f5a660;
    ram_cell[     571] = 32'h4ad10ca8;
    ram_cell[     572] = 32'h419eef37;
    ram_cell[     573] = 32'h2354908a;
    ram_cell[     574] = 32'h61c515cd;
    ram_cell[     575] = 32'h7f4ea6a4;
    ram_cell[     576] = 32'h0973effb;
    ram_cell[     577] = 32'he349923a;
    ram_cell[     578] = 32'h44cea500;
    ram_cell[     579] = 32'h97012dfe;
    ram_cell[     580] = 32'h45c52c73;
    ram_cell[     581] = 32'hd2ba1525;
    ram_cell[     582] = 32'h30983689;
    ram_cell[     583] = 32'h26cd2e0e;
    ram_cell[     584] = 32'h4f52af80;
    ram_cell[     585] = 32'h88e11a4b;
    ram_cell[     586] = 32'h25bd245f;
    ram_cell[     587] = 32'h2c5bd0ab;
    ram_cell[     588] = 32'h968e1339;
    ram_cell[     589] = 32'h288dd031;
    ram_cell[     590] = 32'h0b9df549;
    ram_cell[     591] = 32'h433750e9;
    ram_cell[     592] = 32'h266a6969;
    ram_cell[     593] = 32'h52f6cb76;
    ram_cell[     594] = 32'ha8420dee;
    ram_cell[     595] = 32'h72d12cf5;
    ram_cell[     596] = 32'h61a05b12;
    ram_cell[     597] = 32'hd8468da8;
    ram_cell[     598] = 32'h5a435b49;
    ram_cell[     599] = 32'hff321543;
    ram_cell[     600] = 32'h12d93243;
    ram_cell[     601] = 32'h845a0341;
    ram_cell[     602] = 32'h3517b214;
    ram_cell[     603] = 32'h1c088092;
    ram_cell[     604] = 32'h2394c980;
    ram_cell[     605] = 32'hf3e54683;
    ram_cell[     606] = 32'h05d457e3;
    ram_cell[     607] = 32'h33100d0a;
    ram_cell[     608] = 32'hd2a651d0;
    ram_cell[     609] = 32'hf9eea12c;
    ram_cell[     610] = 32'h484d0459;
    ram_cell[     611] = 32'h4b06a223;
    ram_cell[     612] = 32'he7ab4133;
    ram_cell[     613] = 32'h3054eced;
    ram_cell[     614] = 32'h89cd5106;
    ram_cell[     615] = 32'h66b6ed93;
    ram_cell[     616] = 32'h7227dbcc;
    ram_cell[     617] = 32'h5b20cfe9;
    ram_cell[     618] = 32'hca3da191;
    ram_cell[     619] = 32'hd3edef06;
    ram_cell[     620] = 32'h715206fd;
    ram_cell[     621] = 32'h0e84785b;
    ram_cell[     622] = 32'h6bf10b8e;
    ram_cell[     623] = 32'h839b9356;
    ram_cell[     624] = 32'hb94c0165;
    ram_cell[     625] = 32'h423b8d13;
    ram_cell[     626] = 32'h8060d6dd;
    ram_cell[     627] = 32'hff9c5a4a;
    ram_cell[     628] = 32'h53840267;
    ram_cell[     629] = 32'h431691c6;
    ram_cell[     630] = 32'hafc9ca71;
    ram_cell[     631] = 32'h72af66b8;
    ram_cell[     632] = 32'h54e53b40;
    ram_cell[     633] = 32'h2453d718;
    ram_cell[     634] = 32'h9d8ed9db;
    ram_cell[     635] = 32'h22cb669e;
    ram_cell[     636] = 32'h25495e11;
    ram_cell[     637] = 32'hb2cd618a;
    ram_cell[     638] = 32'h5a4d0242;
    ram_cell[     639] = 32'h3bc06731;
    ram_cell[     640] = 32'h0022aebd;
    ram_cell[     641] = 32'hd7d8344c;
    ram_cell[     642] = 32'hbb11596c;
    ram_cell[     643] = 32'h6476bf8c;
    ram_cell[     644] = 32'hf5e69587;
    ram_cell[     645] = 32'h1460f4f7;
    ram_cell[     646] = 32'h78ad0740;
    ram_cell[     647] = 32'hcf6e2f54;
    ram_cell[     648] = 32'h0987fa21;
    ram_cell[     649] = 32'h6bfda3b7;
    ram_cell[     650] = 32'h56d4b30e;
    ram_cell[     651] = 32'h2a158757;
    ram_cell[     652] = 32'h0f76c8e0;
    ram_cell[     653] = 32'hd7adbec5;
    ram_cell[     654] = 32'ha97f732e;
    ram_cell[     655] = 32'h8b11a7d3;
    ram_cell[     656] = 32'h0fb5f10c;
    ram_cell[     657] = 32'h5ba1a1df;
    ram_cell[     658] = 32'h90a31b34;
    ram_cell[     659] = 32'h44001ea3;
    ram_cell[     660] = 32'heb63947f;
    ram_cell[     661] = 32'heac97cc1;
    ram_cell[     662] = 32'h30e220f8;
    ram_cell[     663] = 32'hd7d46a95;
    ram_cell[     664] = 32'h224d1c17;
    ram_cell[     665] = 32'h8a8fb287;
    ram_cell[     666] = 32'hf31e9f8e;
    ram_cell[     667] = 32'hf35cbb08;
    ram_cell[     668] = 32'he42e9e26;
    ram_cell[     669] = 32'hd7cb6a8e;
    ram_cell[     670] = 32'h5b906db0;
    ram_cell[     671] = 32'hf973461b;
    ram_cell[     672] = 32'he112049b;
    ram_cell[     673] = 32'hd99d65ed;
    ram_cell[     674] = 32'hced25155;
    ram_cell[     675] = 32'h28c4a308;
    ram_cell[     676] = 32'h286b92f9;
    ram_cell[     677] = 32'he502f2f6;
    ram_cell[     678] = 32'h02d8b83e;
    ram_cell[     679] = 32'h60d50190;
    ram_cell[     680] = 32'ha9de21c2;
    ram_cell[     681] = 32'h404f2082;
    ram_cell[     682] = 32'heaca49c4;
    ram_cell[     683] = 32'hb113730a;
    ram_cell[     684] = 32'hcd938f53;
    ram_cell[     685] = 32'h507d3f3c;
    ram_cell[     686] = 32'hd9eb4caa;
    ram_cell[     687] = 32'hfccbd727;
    ram_cell[     688] = 32'h6fbcf5d8;
    ram_cell[     689] = 32'hefed9797;
    ram_cell[     690] = 32'he5346e43;
    ram_cell[     691] = 32'h76113d25;
    ram_cell[     692] = 32'h8e7868d8;
    ram_cell[     693] = 32'h5aeb5b07;
    ram_cell[     694] = 32'h664fdb51;
    ram_cell[     695] = 32'hb1223fff;
    ram_cell[     696] = 32'h4a4c12c9;
    ram_cell[     697] = 32'h02ca1830;
    ram_cell[     698] = 32'h081240a7;
    ram_cell[     699] = 32'h45ff2c86;
    ram_cell[     700] = 32'hce8970fd;
    ram_cell[     701] = 32'h391ba364;
    ram_cell[     702] = 32'h87a95ee6;
    ram_cell[     703] = 32'h6e4b050c;
    ram_cell[     704] = 32'hc1802273;
    ram_cell[     705] = 32'h9cd5d25e;
    ram_cell[     706] = 32'hde97e3e9;
    ram_cell[     707] = 32'hc28bcbd8;
    ram_cell[     708] = 32'h87c2700b;
    ram_cell[     709] = 32'h5e1a6292;
    ram_cell[     710] = 32'h165b312c;
    ram_cell[     711] = 32'hb7e1be03;
    ram_cell[     712] = 32'heffc520a;
    ram_cell[     713] = 32'hbf7cb747;
    ram_cell[     714] = 32'hf2180965;
    ram_cell[     715] = 32'hb22a44c0;
    ram_cell[     716] = 32'h074dc273;
    ram_cell[     717] = 32'hf09188be;
    ram_cell[     718] = 32'h07498d3d;
    ram_cell[     719] = 32'hfaf98376;
    ram_cell[     720] = 32'h5da42487;
    ram_cell[     721] = 32'hc0507427;
    ram_cell[     722] = 32'h6d552e6c;
    ram_cell[     723] = 32'h2518eca5;
    ram_cell[     724] = 32'hdee2e7c2;
    ram_cell[     725] = 32'h08103049;
    ram_cell[     726] = 32'hc1acf0c7;
    ram_cell[     727] = 32'h86c15151;
    ram_cell[     728] = 32'hec4ec34b;
    ram_cell[     729] = 32'h1e592dad;
    ram_cell[     730] = 32'h548aa690;
    ram_cell[     731] = 32'h26cfeb40;
    ram_cell[     732] = 32'h4abb6035;
    ram_cell[     733] = 32'hf3e6f84f;
    ram_cell[     734] = 32'hb96d6262;
    ram_cell[     735] = 32'h88038fc0;
    ram_cell[     736] = 32'h048e097b;
    ram_cell[     737] = 32'h5fabad33;
    ram_cell[     738] = 32'he1866c0d;
    ram_cell[     739] = 32'hc6a820fb;
    ram_cell[     740] = 32'hacaf2536;
    ram_cell[     741] = 32'h9e5af517;
    ram_cell[     742] = 32'h8562638e;
    ram_cell[     743] = 32'hfe74798f;
    ram_cell[     744] = 32'hdd8f11aa;
    ram_cell[     745] = 32'h45dab01b;
    ram_cell[     746] = 32'heec1103f;
    ram_cell[     747] = 32'h6fb1b9f7;
    ram_cell[     748] = 32'he4cddf91;
    ram_cell[     749] = 32'h79dcf2d4;
    ram_cell[     750] = 32'h17f36be4;
    ram_cell[     751] = 32'h3da80dfb;
    ram_cell[     752] = 32'h6794f5a1;
    ram_cell[     753] = 32'he68f8669;
    ram_cell[     754] = 32'h4f1410c5;
    ram_cell[     755] = 32'h12c79cd7;
    ram_cell[     756] = 32'hb667c3f2;
    ram_cell[     757] = 32'h6d440d26;
    ram_cell[     758] = 32'h8fd07707;
    ram_cell[     759] = 32'ha76a310d;
    ram_cell[     760] = 32'heeccf41c;
    ram_cell[     761] = 32'h08f4c4eb;
    ram_cell[     762] = 32'h58cff8f2;
    ram_cell[     763] = 32'h4f7af8b7;
    ram_cell[     764] = 32'h5906fb04;
    ram_cell[     765] = 32'h8b7d88a0;
    ram_cell[     766] = 32'hd2f3fbf8;
    ram_cell[     767] = 32'h3dfdd8b0;
end

endmodule

