
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h2d0f83ed;
    ram_cell[       1] = 32'h0;  // 32'h33a87d57;
    ram_cell[       2] = 32'h0;  // 32'h5d31eb66;
    ram_cell[       3] = 32'h0;  // 32'h003408e3;
    ram_cell[       4] = 32'h0;  // 32'h27e711c0;
    ram_cell[       5] = 32'h0;  // 32'h5904d6f3;
    ram_cell[       6] = 32'h0;  // 32'h161c0157;
    ram_cell[       7] = 32'h0;  // 32'h5696304e;
    ram_cell[       8] = 32'h0;  // 32'h0f607ac0;
    ram_cell[       9] = 32'h0;  // 32'h17b5c6c6;
    ram_cell[      10] = 32'h0;  // 32'hfb4fbb3d;
    ram_cell[      11] = 32'h0;  // 32'hb084071e;
    ram_cell[      12] = 32'h0;  // 32'h72c537a1;
    ram_cell[      13] = 32'h0;  // 32'hb02f196d;
    ram_cell[      14] = 32'h0;  // 32'h4b10b345;
    ram_cell[      15] = 32'h0;  // 32'had34c0e3;
    ram_cell[      16] = 32'h0;  // 32'hbb065aaa;
    ram_cell[      17] = 32'h0;  // 32'h23c4972c;
    ram_cell[      18] = 32'h0;  // 32'h2e2033dd;
    ram_cell[      19] = 32'h0;  // 32'h2d894445;
    ram_cell[      20] = 32'h0;  // 32'h1088bc9f;
    ram_cell[      21] = 32'h0;  // 32'h375b46c0;
    ram_cell[      22] = 32'h0;  // 32'ha48b9beb;
    ram_cell[      23] = 32'h0;  // 32'h6eaf54c0;
    ram_cell[      24] = 32'h0;  // 32'he821dcae;
    ram_cell[      25] = 32'h0;  // 32'h4b5707e1;
    ram_cell[      26] = 32'h0;  // 32'h1ef0cb84;
    ram_cell[      27] = 32'h0;  // 32'hcc598346;
    ram_cell[      28] = 32'h0;  // 32'h1f5aa58d;
    ram_cell[      29] = 32'h0;  // 32'h6de8a783;
    ram_cell[      30] = 32'h0;  // 32'h8506c0b8;
    ram_cell[      31] = 32'h0;  // 32'h7d877571;
    ram_cell[      32] = 32'h0;  // 32'h4f1475e6;
    ram_cell[      33] = 32'h0;  // 32'hc73b269c;
    ram_cell[      34] = 32'h0;  // 32'h89efa412;
    ram_cell[      35] = 32'h0;  // 32'haf30f84d;
    ram_cell[      36] = 32'h0;  // 32'hf6c4cb06;
    ram_cell[      37] = 32'h0;  // 32'he547d90b;
    ram_cell[      38] = 32'h0;  // 32'hfce21254;
    ram_cell[      39] = 32'h0;  // 32'h3050f925;
    ram_cell[      40] = 32'h0;  // 32'hf7c2a797;
    ram_cell[      41] = 32'h0;  // 32'hdb4cffba;
    ram_cell[      42] = 32'h0;  // 32'h6796d1b4;
    ram_cell[      43] = 32'h0;  // 32'h41c231aa;
    ram_cell[      44] = 32'h0;  // 32'h9b90179e;
    ram_cell[      45] = 32'h0;  // 32'h2cc2cb2e;
    ram_cell[      46] = 32'h0;  // 32'hace5a079;
    ram_cell[      47] = 32'h0;  // 32'h64e15f6b;
    ram_cell[      48] = 32'h0;  // 32'h3a8ea522;
    ram_cell[      49] = 32'h0;  // 32'h1f842b28;
    ram_cell[      50] = 32'h0;  // 32'hebd85223;
    ram_cell[      51] = 32'h0;  // 32'hf55b200d;
    ram_cell[      52] = 32'h0;  // 32'hd1eb11b6;
    ram_cell[      53] = 32'h0;  // 32'hd249d662;
    ram_cell[      54] = 32'h0;  // 32'h68eee00b;
    ram_cell[      55] = 32'h0;  // 32'h7398ad54;
    ram_cell[      56] = 32'h0;  // 32'h1a02a837;
    ram_cell[      57] = 32'h0;  // 32'h36aeeebb;
    ram_cell[      58] = 32'h0;  // 32'h1d36f610;
    ram_cell[      59] = 32'h0;  // 32'h4038a555;
    ram_cell[      60] = 32'h0;  // 32'h7dbf7f40;
    ram_cell[      61] = 32'h0;  // 32'h235c327f;
    ram_cell[      62] = 32'h0;  // 32'h81d323d1;
    ram_cell[      63] = 32'h0;  // 32'hd74a47db;
    ram_cell[      64] = 32'h0;  // 32'hd0ec8a1e;
    ram_cell[      65] = 32'h0;  // 32'hb4dfe7ec;
    ram_cell[      66] = 32'h0;  // 32'ha2b90545;
    ram_cell[      67] = 32'h0;  // 32'h763016fa;
    ram_cell[      68] = 32'h0;  // 32'h8a1416f1;
    ram_cell[      69] = 32'h0;  // 32'hffd1762f;
    ram_cell[      70] = 32'h0;  // 32'h731374c1;
    ram_cell[      71] = 32'h0;  // 32'h27e018d2;
    ram_cell[      72] = 32'h0;  // 32'h697c6dea;
    ram_cell[      73] = 32'h0;  // 32'h32b55820;
    ram_cell[      74] = 32'h0;  // 32'he523a953;
    ram_cell[      75] = 32'h0;  // 32'h5ece4621;
    ram_cell[      76] = 32'h0;  // 32'h7c01150b;
    ram_cell[      77] = 32'h0;  // 32'hf8208cad;
    ram_cell[      78] = 32'h0;  // 32'hc656de29;
    ram_cell[      79] = 32'h0;  // 32'h8ba34707;
    ram_cell[      80] = 32'h0;  // 32'hac6873f1;
    ram_cell[      81] = 32'h0;  // 32'hc23eecc9;
    ram_cell[      82] = 32'h0;  // 32'h08fb99ff;
    ram_cell[      83] = 32'h0;  // 32'h959470a5;
    ram_cell[      84] = 32'h0;  // 32'h1fcaf10b;
    ram_cell[      85] = 32'h0;  // 32'h1ae9e95a;
    ram_cell[      86] = 32'h0;  // 32'had48a4be;
    ram_cell[      87] = 32'h0;  // 32'hace88325;
    ram_cell[      88] = 32'h0;  // 32'hed792f4b;
    ram_cell[      89] = 32'h0;  // 32'h9ec76db8;
    ram_cell[      90] = 32'h0;  // 32'h6862f981;
    ram_cell[      91] = 32'h0;  // 32'hc2e3ff54;
    ram_cell[      92] = 32'h0;  // 32'h42b2bdba;
    ram_cell[      93] = 32'h0;  // 32'h14e5264b;
    ram_cell[      94] = 32'h0;  // 32'h91c651e7;
    ram_cell[      95] = 32'h0;  // 32'h6ac8ab0a;
    ram_cell[      96] = 32'h0;  // 32'h2c787282;
    ram_cell[      97] = 32'h0;  // 32'he1aabcba;
    ram_cell[      98] = 32'h0;  // 32'he5aa838c;
    ram_cell[      99] = 32'h0;  // 32'hd6c423c5;
    ram_cell[     100] = 32'h0;  // 32'hcba85f2f;
    ram_cell[     101] = 32'h0;  // 32'hb78ef5e1;
    ram_cell[     102] = 32'h0;  // 32'h0f1775e7;
    ram_cell[     103] = 32'h0;  // 32'hd35d4e47;
    ram_cell[     104] = 32'h0;  // 32'hb8f8eeed;
    ram_cell[     105] = 32'h0;  // 32'ha834d5ca;
    ram_cell[     106] = 32'h0;  // 32'h012c4a1b;
    ram_cell[     107] = 32'h0;  // 32'h3eb77178;
    ram_cell[     108] = 32'h0;  // 32'h69f4a369;
    ram_cell[     109] = 32'h0;  // 32'hd3539dc5;
    ram_cell[     110] = 32'h0;  // 32'h877053d6;
    ram_cell[     111] = 32'h0;  // 32'h56683ca1;
    ram_cell[     112] = 32'h0;  // 32'h684a622b;
    ram_cell[     113] = 32'h0;  // 32'h7e1b778d;
    ram_cell[     114] = 32'h0;  // 32'heb6e6c7b;
    ram_cell[     115] = 32'h0;  // 32'h27b24284;
    ram_cell[     116] = 32'h0;  // 32'h2a93389b;
    ram_cell[     117] = 32'h0;  // 32'h26024649;
    ram_cell[     118] = 32'h0;  // 32'he17f72cb;
    ram_cell[     119] = 32'h0;  // 32'h98e61501;
    ram_cell[     120] = 32'h0;  // 32'h90066125;
    ram_cell[     121] = 32'h0;  // 32'h3cebccf5;
    ram_cell[     122] = 32'h0;  // 32'h3e3d575c;
    ram_cell[     123] = 32'h0;  // 32'ha08efcb7;
    ram_cell[     124] = 32'h0;  // 32'hea8e18ee;
    ram_cell[     125] = 32'h0;  // 32'h27b6a935;
    ram_cell[     126] = 32'h0;  // 32'hf99cf36b;
    ram_cell[     127] = 32'h0;  // 32'h1a3d86b8;
    ram_cell[     128] = 32'h0;  // 32'ha2c26512;
    ram_cell[     129] = 32'h0;  // 32'h41e47f9e;
    ram_cell[     130] = 32'h0;  // 32'h83d16377;
    ram_cell[     131] = 32'h0;  // 32'h409ca205;
    ram_cell[     132] = 32'h0;  // 32'hdcd12bad;
    ram_cell[     133] = 32'h0;  // 32'h175d7b0a;
    ram_cell[     134] = 32'h0;  // 32'h54e99538;
    ram_cell[     135] = 32'h0;  // 32'hb6aa4949;
    ram_cell[     136] = 32'h0;  // 32'h34e357a3;
    ram_cell[     137] = 32'h0;  // 32'hf45cd5c3;
    ram_cell[     138] = 32'h0;  // 32'hefd07754;
    ram_cell[     139] = 32'h0;  // 32'h2cc19b8b;
    ram_cell[     140] = 32'h0;  // 32'h38655607;
    ram_cell[     141] = 32'h0;  // 32'h9cdcdf29;
    ram_cell[     142] = 32'h0;  // 32'h9ccb7347;
    ram_cell[     143] = 32'h0;  // 32'he780972f;
    ram_cell[     144] = 32'h0;  // 32'h7d3d90d2;
    ram_cell[     145] = 32'h0;  // 32'h71efc2d3;
    ram_cell[     146] = 32'h0;  // 32'hd38a6701;
    ram_cell[     147] = 32'h0;  // 32'h6f4175d9;
    ram_cell[     148] = 32'h0;  // 32'h6ff2b2e9;
    ram_cell[     149] = 32'h0;  // 32'h1de995c6;
    ram_cell[     150] = 32'h0;  // 32'hfa05a117;
    ram_cell[     151] = 32'h0;  // 32'h733adfb9;
    ram_cell[     152] = 32'h0;  // 32'h04126623;
    ram_cell[     153] = 32'h0;  // 32'h5cae6e53;
    ram_cell[     154] = 32'h0;  // 32'h19970d72;
    ram_cell[     155] = 32'h0;  // 32'h9a8884bd;
    ram_cell[     156] = 32'h0;  // 32'hf1a96681;
    ram_cell[     157] = 32'h0;  // 32'h6caefcce;
    ram_cell[     158] = 32'h0;  // 32'h5b166e06;
    ram_cell[     159] = 32'h0;  // 32'hf5bfb042;
    ram_cell[     160] = 32'h0;  // 32'hc8ee9c65;
    ram_cell[     161] = 32'h0;  // 32'h972630b9;
    ram_cell[     162] = 32'h0;  // 32'hb476039e;
    ram_cell[     163] = 32'h0;  // 32'h7d3c99b8;
    ram_cell[     164] = 32'h0;  // 32'h56b320b4;
    ram_cell[     165] = 32'h0;  // 32'hdc491f76;
    ram_cell[     166] = 32'h0;  // 32'had290cf7;
    ram_cell[     167] = 32'h0;  // 32'hf795c90a;
    ram_cell[     168] = 32'h0;  // 32'h163edc53;
    ram_cell[     169] = 32'h0;  // 32'h22881f24;
    ram_cell[     170] = 32'h0;  // 32'h9990ec26;
    ram_cell[     171] = 32'h0;  // 32'hb21fb25f;
    ram_cell[     172] = 32'h0;  // 32'h27f6b88f;
    ram_cell[     173] = 32'h0;  // 32'hbc7ff90e;
    ram_cell[     174] = 32'h0;  // 32'h4310d712;
    ram_cell[     175] = 32'h0;  // 32'hfc6d88b3;
    ram_cell[     176] = 32'h0;  // 32'hc04c0cf3;
    ram_cell[     177] = 32'h0;  // 32'hbf031c0e;
    ram_cell[     178] = 32'h0;  // 32'hf83430c1;
    ram_cell[     179] = 32'h0;  // 32'h034df4a2;
    ram_cell[     180] = 32'h0;  // 32'h729d92b0;
    ram_cell[     181] = 32'h0;  // 32'h354406c1;
    ram_cell[     182] = 32'h0;  // 32'h142f35a6;
    ram_cell[     183] = 32'h0;  // 32'h73ee617a;
    ram_cell[     184] = 32'h0;  // 32'h8c259436;
    ram_cell[     185] = 32'h0;  // 32'h1d604b24;
    ram_cell[     186] = 32'h0;  // 32'hd0d3ed7f;
    ram_cell[     187] = 32'h0;  // 32'h2a80bd7c;
    ram_cell[     188] = 32'h0;  // 32'h5104b5ec;
    ram_cell[     189] = 32'h0;  // 32'h3b52e922;
    ram_cell[     190] = 32'h0;  // 32'ha9c542de;
    ram_cell[     191] = 32'h0;  // 32'h995feb18;
    ram_cell[     192] = 32'h0;  // 32'hc7dcca50;
    ram_cell[     193] = 32'h0;  // 32'h65ad6981;
    ram_cell[     194] = 32'h0;  // 32'hf8cade91;
    ram_cell[     195] = 32'h0;  // 32'h6ceef637;
    ram_cell[     196] = 32'h0;  // 32'hbfc04579;
    ram_cell[     197] = 32'h0;  // 32'hd34efaa6;
    ram_cell[     198] = 32'h0;  // 32'h7d2b3e44;
    ram_cell[     199] = 32'h0;  // 32'he9a231f2;
    ram_cell[     200] = 32'h0;  // 32'ha6c2e5af;
    ram_cell[     201] = 32'h0;  // 32'h2e04d979;
    ram_cell[     202] = 32'h0;  // 32'hf9b6e993;
    ram_cell[     203] = 32'h0;  // 32'hea439e62;
    ram_cell[     204] = 32'h0;  // 32'h0ea47e3a;
    ram_cell[     205] = 32'h0;  // 32'hbc58b132;
    ram_cell[     206] = 32'h0;  // 32'ha2e35082;
    ram_cell[     207] = 32'h0;  // 32'h26896313;
    ram_cell[     208] = 32'h0;  // 32'h7df7e380;
    ram_cell[     209] = 32'h0;  // 32'ha688c0fc;
    ram_cell[     210] = 32'h0;  // 32'hea4968c7;
    ram_cell[     211] = 32'h0;  // 32'hbbbc5314;
    ram_cell[     212] = 32'h0;  // 32'hb4678ee2;
    ram_cell[     213] = 32'h0;  // 32'h9fb20234;
    ram_cell[     214] = 32'h0;  // 32'h9b41c3b8;
    ram_cell[     215] = 32'h0;  // 32'h77e8b04c;
    ram_cell[     216] = 32'h0;  // 32'h75401af5;
    ram_cell[     217] = 32'h0;  // 32'hb62666a0;
    ram_cell[     218] = 32'h0;  // 32'h9f6e730e;
    ram_cell[     219] = 32'h0;  // 32'h4d0d8fc9;
    ram_cell[     220] = 32'h0;  // 32'he9306910;
    ram_cell[     221] = 32'h0;  // 32'hea579427;
    ram_cell[     222] = 32'h0;  // 32'hef4e2c89;
    ram_cell[     223] = 32'h0;  // 32'h05773317;
    ram_cell[     224] = 32'h0;  // 32'hc7f04e12;
    ram_cell[     225] = 32'h0;  // 32'h301aea2c;
    ram_cell[     226] = 32'h0;  // 32'h7706579a;
    ram_cell[     227] = 32'h0;  // 32'hfc8e484e;
    ram_cell[     228] = 32'h0;  // 32'h3ef87fe0;
    ram_cell[     229] = 32'h0;  // 32'h034c033d;
    ram_cell[     230] = 32'h0;  // 32'h9567b1b1;
    ram_cell[     231] = 32'h0;  // 32'h0021153b;
    ram_cell[     232] = 32'h0;  // 32'haa8089ba;
    ram_cell[     233] = 32'h0;  // 32'hb0dc51e2;
    ram_cell[     234] = 32'h0;  // 32'he018114f;
    ram_cell[     235] = 32'h0;  // 32'h6134ed56;
    ram_cell[     236] = 32'h0;  // 32'hf2aaec6a;
    ram_cell[     237] = 32'h0;  // 32'h8aca99bf;
    ram_cell[     238] = 32'h0;  // 32'hfa3d9622;
    ram_cell[     239] = 32'h0;  // 32'heec83bd9;
    ram_cell[     240] = 32'h0;  // 32'h17b4128c;
    ram_cell[     241] = 32'h0;  // 32'had97d155;
    ram_cell[     242] = 32'h0;  // 32'hea4d8979;
    ram_cell[     243] = 32'h0;  // 32'h5302a8d2;
    ram_cell[     244] = 32'h0;  // 32'h330ee1f0;
    ram_cell[     245] = 32'h0;  // 32'h2d84a7c0;
    ram_cell[     246] = 32'h0;  // 32'he63023f1;
    ram_cell[     247] = 32'h0;  // 32'ha6045a32;
    ram_cell[     248] = 32'h0;  // 32'h5c8dca96;
    ram_cell[     249] = 32'h0;  // 32'h790be99b;
    ram_cell[     250] = 32'h0;  // 32'h218bdff3;
    ram_cell[     251] = 32'h0;  // 32'h1fed4cdf;
    ram_cell[     252] = 32'h0;  // 32'h99de58c0;
    ram_cell[     253] = 32'h0;  // 32'h7133efc0;
    ram_cell[     254] = 32'h0;  // 32'h5764b036;
    ram_cell[     255] = 32'h0;  // 32'hb1c97f0b;
    // src matrix A
    ram_cell[     256] = 32'hfe5ce7ec;
    ram_cell[     257] = 32'h7c616c7c;
    ram_cell[     258] = 32'h667dad85;
    ram_cell[     259] = 32'hf7444dda;
    ram_cell[     260] = 32'hd8a3eb3a;
    ram_cell[     261] = 32'hc9058ac8;
    ram_cell[     262] = 32'hd0256ee3;
    ram_cell[     263] = 32'h66bf76fc;
    ram_cell[     264] = 32'h7a638176;
    ram_cell[     265] = 32'h74d4e712;
    ram_cell[     266] = 32'h0901c087;
    ram_cell[     267] = 32'h30a242d6;
    ram_cell[     268] = 32'hc2bcc002;
    ram_cell[     269] = 32'h5ceca12b;
    ram_cell[     270] = 32'hc5b535da;
    ram_cell[     271] = 32'h7270b53a;
    ram_cell[     272] = 32'h033d3b5a;
    ram_cell[     273] = 32'h7141bc25;
    ram_cell[     274] = 32'h12a126bb;
    ram_cell[     275] = 32'hba124757;
    ram_cell[     276] = 32'hc7b31163;
    ram_cell[     277] = 32'h21a299ce;
    ram_cell[     278] = 32'ha5f14601;
    ram_cell[     279] = 32'hc4d99442;
    ram_cell[     280] = 32'h1b2c3380;
    ram_cell[     281] = 32'h20f3ee4a;
    ram_cell[     282] = 32'ha11e017b;
    ram_cell[     283] = 32'h94cdec9a;
    ram_cell[     284] = 32'he4dd6907;
    ram_cell[     285] = 32'hdc7ef635;
    ram_cell[     286] = 32'h7518058c;
    ram_cell[     287] = 32'h4ed20093;
    ram_cell[     288] = 32'h28a6940e;
    ram_cell[     289] = 32'h6a8617bf;
    ram_cell[     290] = 32'h068b08e0;
    ram_cell[     291] = 32'h5876d8f9;
    ram_cell[     292] = 32'h09ee1237;
    ram_cell[     293] = 32'hc9258ad5;
    ram_cell[     294] = 32'h059203de;
    ram_cell[     295] = 32'hb3744ada;
    ram_cell[     296] = 32'h67bf111c;
    ram_cell[     297] = 32'h9efe4acf;
    ram_cell[     298] = 32'ha901e544;
    ram_cell[     299] = 32'h303c7f16;
    ram_cell[     300] = 32'ha5aae4cc;
    ram_cell[     301] = 32'hb0635bcd;
    ram_cell[     302] = 32'he7579159;
    ram_cell[     303] = 32'h18ec40ae;
    ram_cell[     304] = 32'hed42907f;
    ram_cell[     305] = 32'h9684dce8;
    ram_cell[     306] = 32'hae5ce088;
    ram_cell[     307] = 32'ha312bca4;
    ram_cell[     308] = 32'h9595878c;
    ram_cell[     309] = 32'h89409011;
    ram_cell[     310] = 32'h09cf0951;
    ram_cell[     311] = 32'hda2c449d;
    ram_cell[     312] = 32'hcdc852a9;
    ram_cell[     313] = 32'hdf2d369e;
    ram_cell[     314] = 32'h262db29a;
    ram_cell[     315] = 32'h0d3326e9;
    ram_cell[     316] = 32'h0d062e06;
    ram_cell[     317] = 32'hae7c41bd;
    ram_cell[     318] = 32'h5fa453b4;
    ram_cell[     319] = 32'hb3f2b170;
    ram_cell[     320] = 32'h725780b4;
    ram_cell[     321] = 32'hf6e1192b;
    ram_cell[     322] = 32'h124f393a;
    ram_cell[     323] = 32'h1ef8d079;
    ram_cell[     324] = 32'he2c0d1f5;
    ram_cell[     325] = 32'hb6823aae;
    ram_cell[     326] = 32'h386e62f4;
    ram_cell[     327] = 32'hd0db0211;
    ram_cell[     328] = 32'h94351946;
    ram_cell[     329] = 32'he949d429;
    ram_cell[     330] = 32'h5a8e2158;
    ram_cell[     331] = 32'h810f4488;
    ram_cell[     332] = 32'h644a2590;
    ram_cell[     333] = 32'h82d2d0f1;
    ram_cell[     334] = 32'h0c2e0bc4;
    ram_cell[     335] = 32'h23a0f68b;
    ram_cell[     336] = 32'h1071d666;
    ram_cell[     337] = 32'h3ab280ec;
    ram_cell[     338] = 32'h34f79102;
    ram_cell[     339] = 32'hf461d141;
    ram_cell[     340] = 32'hb3f551e0;
    ram_cell[     341] = 32'h1e033fd7;
    ram_cell[     342] = 32'h78ffa5b5;
    ram_cell[     343] = 32'hb2be2b73;
    ram_cell[     344] = 32'h69aaa948;
    ram_cell[     345] = 32'h43d04958;
    ram_cell[     346] = 32'h5b0b3b48;
    ram_cell[     347] = 32'h68327ac5;
    ram_cell[     348] = 32'h5c8cd082;
    ram_cell[     349] = 32'hc67cc4f0;
    ram_cell[     350] = 32'h1c07ea91;
    ram_cell[     351] = 32'hf805c826;
    ram_cell[     352] = 32'h92951893;
    ram_cell[     353] = 32'h68fdd827;
    ram_cell[     354] = 32'ha94ec103;
    ram_cell[     355] = 32'h8fd5f013;
    ram_cell[     356] = 32'h170ef61a;
    ram_cell[     357] = 32'hf7afd767;
    ram_cell[     358] = 32'hd6fa8b84;
    ram_cell[     359] = 32'hdd25b5cf;
    ram_cell[     360] = 32'h3e643e6f;
    ram_cell[     361] = 32'h889d4cc8;
    ram_cell[     362] = 32'habca5a85;
    ram_cell[     363] = 32'h8032f63e;
    ram_cell[     364] = 32'h5babbd32;
    ram_cell[     365] = 32'ha11a3b65;
    ram_cell[     366] = 32'h164dd7ec;
    ram_cell[     367] = 32'hfac09ca5;
    ram_cell[     368] = 32'h4282b933;
    ram_cell[     369] = 32'h4122e01f;
    ram_cell[     370] = 32'h54b2c69e;
    ram_cell[     371] = 32'h3d3dc5e1;
    ram_cell[     372] = 32'h32afc1d3;
    ram_cell[     373] = 32'hbeaecd73;
    ram_cell[     374] = 32'h92c3c142;
    ram_cell[     375] = 32'hfc3a1957;
    ram_cell[     376] = 32'h88cdd8a8;
    ram_cell[     377] = 32'h65512ca7;
    ram_cell[     378] = 32'hfa81f598;
    ram_cell[     379] = 32'hf1897b30;
    ram_cell[     380] = 32'hdcbe0c3d;
    ram_cell[     381] = 32'hdf103fba;
    ram_cell[     382] = 32'h6fc44f52;
    ram_cell[     383] = 32'h232cc768;
    ram_cell[     384] = 32'hebffe3fd;
    ram_cell[     385] = 32'h1276dd42;
    ram_cell[     386] = 32'hc68beb05;
    ram_cell[     387] = 32'h5c9bcc8b;
    ram_cell[     388] = 32'h779069ca;
    ram_cell[     389] = 32'h28ba9c93;
    ram_cell[     390] = 32'h30f791f6;
    ram_cell[     391] = 32'he44db06d;
    ram_cell[     392] = 32'haea3b461;
    ram_cell[     393] = 32'h17a899d5;
    ram_cell[     394] = 32'h897b29a0;
    ram_cell[     395] = 32'h7b1f11ff;
    ram_cell[     396] = 32'h237d2238;
    ram_cell[     397] = 32'hef9c8bef;
    ram_cell[     398] = 32'he1a5d5b3;
    ram_cell[     399] = 32'hd2ad867c;
    ram_cell[     400] = 32'h9707f323;
    ram_cell[     401] = 32'h27072e23;
    ram_cell[     402] = 32'hbc64e074;
    ram_cell[     403] = 32'ha7020175;
    ram_cell[     404] = 32'hd2301d12;
    ram_cell[     405] = 32'h94e59c56;
    ram_cell[     406] = 32'h251b5f29;
    ram_cell[     407] = 32'h4e8034da;
    ram_cell[     408] = 32'h0ad7dbbf;
    ram_cell[     409] = 32'h3251d26d;
    ram_cell[     410] = 32'h3b63e9c3;
    ram_cell[     411] = 32'h43c0c88d;
    ram_cell[     412] = 32'h03922467;
    ram_cell[     413] = 32'h53351af3;
    ram_cell[     414] = 32'h2996867a;
    ram_cell[     415] = 32'he49df469;
    ram_cell[     416] = 32'h79fc4b57;
    ram_cell[     417] = 32'hea6b18b3;
    ram_cell[     418] = 32'h2e6bff4e;
    ram_cell[     419] = 32'hff491762;
    ram_cell[     420] = 32'h332e4d33;
    ram_cell[     421] = 32'h163d54d2;
    ram_cell[     422] = 32'h09d7a2e5;
    ram_cell[     423] = 32'h703709f0;
    ram_cell[     424] = 32'hba411886;
    ram_cell[     425] = 32'h978bf814;
    ram_cell[     426] = 32'he2912229;
    ram_cell[     427] = 32'h40f92942;
    ram_cell[     428] = 32'h292d7e05;
    ram_cell[     429] = 32'hb0498a35;
    ram_cell[     430] = 32'hececfeeb;
    ram_cell[     431] = 32'hf68bc1b9;
    ram_cell[     432] = 32'h598cf927;
    ram_cell[     433] = 32'h2dc7609a;
    ram_cell[     434] = 32'h55f4d444;
    ram_cell[     435] = 32'h2be173d8;
    ram_cell[     436] = 32'h2e27852f;
    ram_cell[     437] = 32'h851c3f2c;
    ram_cell[     438] = 32'ha815def2;
    ram_cell[     439] = 32'h092e0a80;
    ram_cell[     440] = 32'hc99649ca;
    ram_cell[     441] = 32'h3f517af8;
    ram_cell[     442] = 32'h96383bae;
    ram_cell[     443] = 32'hc489d924;
    ram_cell[     444] = 32'hcec2fd18;
    ram_cell[     445] = 32'h677f5556;
    ram_cell[     446] = 32'h81aacec8;
    ram_cell[     447] = 32'h57502af7;
    ram_cell[     448] = 32'h077657a8;
    ram_cell[     449] = 32'h24f771d8;
    ram_cell[     450] = 32'hf225599a;
    ram_cell[     451] = 32'hb2ce289d;
    ram_cell[     452] = 32'hd19343c4;
    ram_cell[     453] = 32'hf8ee628e;
    ram_cell[     454] = 32'h802c4571;
    ram_cell[     455] = 32'h6e59b61d;
    ram_cell[     456] = 32'h73da9e1f;
    ram_cell[     457] = 32'hc0216758;
    ram_cell[     458] = 32'h063d0e36;
    ram_cell[     459] = 32'he9c20e5b;
    ram_cell[     460] = 32'hd05b4da9;
    ram_cell[     461] = 32'hb46b3571;
    ram_cell[     462] = 32'h747a159e;
    ram_cell[     463] = 32'h84917a96;
    ram_cell[     464] = 32'ha7e5801a;
    ram_cell[     465] = 32'hfbee07ad;
    ram_cell[     466] = 32'h65b3510e;
    ram_cell[     467] = 32'h6d4e8b34;
    ram_cell[     468] = 32'h01130200;
    ram_cell[     469] = 32'hac314907;
    ram_cell[     470] = 32'h25d35368;
    ram_cell[     471] = 32'ha04a48bf;
    ram_cell[     472] = 32'h615d3a55;
    ram_cell[     473] = 32'hc36dfb5f;
    ram_cell[     474] = 32'hadfbf23c;
    ram_cell[     475] = 32'h0e091511;
    ram_cell[     476] = 32'had22541c;
    ram_cell[     477] = 32'heb4b3031;
    ram_cell[     478] = 32'h91c856d9;
    ram_cell[     479] = 32'h9b77d296;
    ram_cell[     480] = 32'h217921be;
    ram_cell[     481] = 32'h167f1f6b;
    ram_cell[     482] = 32'h68b29446;
    ram_cell[     483] = 32'h87c1f4e6;
    ram_cell[     484] = 32'h2a7eb20f;
    ram_cell[     485] = 32'hc3fa2be4;
    ram_cell[     486] = 32'h54b04c38;
    ram_cell[     487] = 32'h42c1f68a;
    ram_cell[     488] = 32'h89029bb3;
    ram_cell[     489] = 32'hdc5fa73a;
    ram_cell[     490] = 32'hd373a596;
    ram_cell[     491] = 32'he3eb6a9c;
    ram_cell[     492] = 32'h342b43b1;
    ram_cell[     493] = 32'hf70dde90;
    ram_cell[     494] = 32'hd5b1f04a;
    ram_cell[     495] = 32'h5e808d97;
    ram_cell[     496] = 32'hc4e10996;
    ram_cell[     497] = 32'h51b7addc;
    ram_cell[     498] = 32'h4e28150d;
    ram_cell[     499] = 32'hdb0f0764;
    ram_cell[     500] = 32'h16b7b15d;
    ram_cell[     501] = 32'h0d92a537;
    ram_cell[     502] = 32'hae9b09c2;
    ram_cell[     503] = 32'h93e6b6cc;
    ram_cell[     504] = 32'h61d69067;
    ram_cell[     505] = 32'hf02206bd;
    ram_cell[     506] = 32'hdc6227f6;
    ram_cell[     507] = 32'hb0635fc0;
    ram_cell[     508] = 32'h92f2c87d;
    ram_cell[     509] = 32'h2e450761;
    ram_cell[     510] = 32'hf3183d5a;
    ram_cell[     511] = 32'he9dff695;
    // src matrix B
    ram_cell[     512] = 32'he97e3c82;
    ram_cell[     513] = 32'hd4950e45;
    ram_cell[     514] = 32'hd70497a2;
    ram_cell[     515] = 32'h40c9ce3a;
    ram_cell[     516] = 32'h6e367c98;
    ram_cell[     517] = 32'hf53698a0;
    ram_cell[     518] = 32'h30cab45e;
    ram_cell[     519] = 32'h340117c6;
    ram_cell[     520] = 32'h14a54292;
    ram_cell[     521] = 32'h14f84120;
    ram_cell[     522] = 32'ha3afa0ff;
    ram_cell[     523] = 32'h246f86b8;
    ram_cell[     524] = 32'h9b3c0951;
    ram_cell[     525] = 32'hf3591958;
    ram_cell[     526] = 32'h2481f987;
    ram_cell[     527] = 32'h431e860a;
    ram_cell[     528] = 32'h39d17803;
    ram_cell[     529] = 32'h27f43810;
    ram_cell[     530] = 32'h447e0f8e;
    ram_cell[     531] = 32'hcc2cf55d;
    ram_cell[     532] = 32'hbebd231c;
    ram_cell[     533] = 32'h213cc1ce;
    ram_cell[     534] = 32'h88d914d7;
    ram_cell[     535] = 32'h2288a242;
    ram_cell[     536] = 32'hddd3727f;
    ram_cell[     537] = 32'h01689ee8;
    ram_cell[     538] = 32'hbb0e737c;
    ram_cell[     539] = 32'h221ea18c;
    ram_cell[     540] = 32'hcaeb7286;
    ram_cell[     541] = 32'h0b832747;
    ram_cell[     542] = 32'ha6de63a3;
    ram_cell[     543] = 32'h4104ce2b;
    ram_cell[     544] = 32'hf52f3ca8;
    ram_cell[     545] = 32'h1b51afbd;
    ram_cell[     546] = 32'h7db84eff;
    ram_cell[     547] = 32'h8a079dc3;
    ram_cell[     548] = 32'h30c92b2b;
    ram_cell[     549] = 32'h032b8f5d;
    ram_cell[     550] = 32'h4e13ecf7;
    ram_cell[     551] = 32'heca57665;
    ram_cell[     552] = 32'h86532888;
    ram_cell[     553] = 32'h087220ba;
    ram_cell[     554] = 32'hab0e8ece;
    ram_cell[     555] = 32'h88392ca9;
    ram_cell[     556] = 32'hcc28e7c7;
    ram_cell[     557] = 32'hb450773b;
    ram_cell[     558] = 32'h4b0d76b1;
    ram_cell[     559] = 32'h2f4412c8;
    ram_cell[     560] = 32'h61241847;
    ram_cell[     561] = 32'hd6486dee;
    ram_cell[     562] = 32'h3e797cff;
    ram_cell[     563] = 32'hf93eb20f;
    ram_cell[     564] = 32'h0c3b3edc;
    ram_cell[     565] = 32'h54411601;
    ram_cell[     566] = 32'h61c4a4f4;
    ram_cell[     567] = 32'h5b9283d0;
    ram_cell[     568] = 32'h16ce9ce9;
    ram_cell[     569] = 32'h001bf4ad;
    ram_cell[     570] = 32'h575a3c03;
    ram_cell[     571] = 32'hd71f6c5b;
    ram_cell[     572] = 32'h5d8a95f7;
    ram_cell[     573] = 32'h2f8c58f4;
    ram_cell[     574] = 32'hf365f111;
    ram_cell[     575] = 32'h8962855f;
    ram_cell[     576] = 32'h93306edb;
    ram_cell[     577] = 32'h1b076835;
    ram_cell[     578] = 32'hc075386c;
    ram_cell[     579] = 32'h328458a4;
    ram_cell[     580] = 32'haaa6120b;
    ram_cell[     581] = 32'h65457450;
    ram_cell[     582] = 32'h9ad5b6d8;
    ram_cell[     583] = 32'h1cdf2550;
    ram_cell[     584] = 32'h87a11ee2;
    ram_cell[     585] = 32'he4b8068c;
    ram_cell[     586] = 32'h2b938bb5;
    ram_cell[     587] = 32'h67d522c0;
    ram_cell[     588] = 32'hf6843941;
    ram_cell[     589] = 32'h57517ca6;
    ram_cell[     590] = 32'h44d17ad0;
    ram_cell[     591] = 32'h4d7f0775;
    ram_cell[     592] = 32'hc743bca1;
    ram_cell[     593] = 32'haceaaaa6;
    ram_cell[     594] = 32'h65438ef2;
    ram_cell[     595] = 32'h5ef69703;
    ram_cell[     596] = 32'h5789b704;
    ram_cell[     597] = 32'h2fa789c6;
    ram_cell[     598] = 32'h477e8428;
    ram_cell[     599] = 32'h8b25c718;
    ram_cell[     600] = 32'h5d6b37ab;
    ram_cell[     601] = 32'h3c0fab29;
    ram_cell[     602] = 32'h08ff9097;
    ram_cell[     603] = 32'h6987685d;
    ram_cell[     604] = 32'hdf9c1070;
    ram_cell[     605] = 32'h940b417c;
    ram_cell[     606] = 32'h2f2fdb5b;
    ram_cell[     607] = 32'h12dad4ed;
    ram_cell[     608] = 32'hd64fda1b;
    ram_cell[     609] = 32'h3a06274a;
    ram_cell[     610] = 32'h4c959c65;
    ram_cell[     611] = 32'h20999ded;
    ram_cell[     612] = 32'h8829cebd;
    ram_cell[     613] = 32'h2b9bf736;
    ram_cell[     614] = 32'hc33d3194;
    ram_cell[     615] = 32'h6b9a53fc;
    ram_cell[     616] = 32'h3e12875d;
    ram_cell[     617] = 32'h507089a7;
    ram_cell[     618] = 32'hc71483ec;
    ram_cell[     619] = 32'h58f26d30;
    ram_cell[     620] = 32'hdfe7bd8d;
    ram_cell[     621] = 32'h3d266cf3;
    ram_cell[     622] = 32'h222d96a7;
    ram_cell[     623] = 32'h394557bf;
    ram_cell[     624] = 32'hdf8cedd3;
    ram_cell[     625] = 32'hc584da11;
    ram_cell[     626] = 32'h0ceb0fc5;
    ram_cell[     627] = 32'h9a749103;
    ram_cell[     628] = 32'h2613fad0;
    ram_cell[     629] = 32'hf5c1a42f;
    ram_cell[     630] = 32'h44e9cf08;
    ram_cell[     631] = 32'he48f1bc0;
    ram_cell[     632] = 32'ha5fdff1c;
    ram_cell[     633] = 32'h1c13d0bd;
    ram_cell[     634] = 32'h97a69be1;
    ram_cell[     635] = 32'h6220de83;
    ram_cell[     636] = 32'h6d3cfea0;
    ram_cell[     637] = 32'h5979abe5;
    ram_cell[     638] = 32'h6aacc249;
    ram_cell[     639] = 32'hfb2da3d7;
    ram_cell[     640] = 32'h5661513a;
    ram_cell[     641] = 32'h3cb4a061;
    ram_cell[     642] = 32'h67532010;
    ram_cell[     643] = 32'h4afae745;
    ram_cell[     644] = 32'h8e02ef0b;
    ram_cell[     645] = 32'h51b280bb;
    ram_cell[     646] = 32'h8599581d;
    ram_cell[     647] = 32'h73b4cac7;
    ram_cell[     648] = 32'hc9ef92d3;
    ram_cell[     649] = 32'hbb280112;
    ram_cell[     650] = 32'h304267e3;
    ram_cell[     651] = 32'h85ff4189;
    ram_cell[     652] = 32'h6bfac6f7;
    ram_cell[     653] = 32'hfcb99cd9;
    ram_cell[     654] = 32'hefac6bde;
    ram_cell[     655] = 32'he419256a;
    ram_cell[     656] = 32'h9cc95aea;
    ram_cell[     657] = 32'h238ab906;
    ram_cell[     658] = 32'ha144309e;
    ram_cell[     659] = 32'h52e94ae4;
    ram_cell[     660] = 32'hdf213d11;
    ram_cell[     661] = 32'h067bdc28;
    ram_cell[     662] = 32'he524f6c1;
    ram_cell[     663] = 32'h2c47fda3;
    ram_cell[     664] = 32'h65f65838;
    ram_cell[     665] = 32'ha2523622;
    ram_cell[     666] = 32'h9477f475;
    ram_cell[     667] = 32'h7e4c4de1;
    ram_cell[     668] = 32'h520653f1;
    ram_cell[     669] = 32'h78e61f16;
    ram_cell[     670] = 32'h0abbfd86;
    ram_cell[     671] = 32'h0c9bcbe5;
    ram_cell[     672] = 32'h224006b0;
    ram_cell[     673] = 32'hdd21a07e;
    ram_cell[     674] = 32'ha5c08c2c;
    ram_cell[     675] = 32'h8ef57674;
    ram_cell[     676] = 32'h62968fa2;
    ram_cell[     677] = 32'h1f5681de;
    ram_cell[     678] = 32'he9386eb9;
    ram_cell[     679] = 32'h45cedad8;
    ram_cell[     680] = 32'hd006eb9d;
    ram_cell[     681] = 32'h993534c7;
    ram_cell[     682] = 32'h293ce67b;
    ram_cell[     683] = 32'h5dda0147;
    ram_cell[     684] = 32'h12ef98cf;
    ram_cell[     685] = 32'hc2692a20;
    ram_cell[     686] = 32'hf4cfd92c;
    ram_cell[     687] = 32'hd5752471;
    ram_cell[     688] = 32'h4ae2e645;
    ram_cell[     689] = 32'he04be703;
    ram_cell[     690] = 32'h95c787e7;
    ram_cell[     691] = 32'h2096154a;
    ram_cell[     692] = 32'h7ad83324;
    ram_cell[     693] = 32'h4b159e16;
    ram_cell[     694] = 32'h6d289bdf;
    ram_cell[     695] = 32'h5103d028;
    ram_cell[     696] = 32'h324c6bc8;
    ram_cell[     697] = 32'h98062052;
    ram_cell[     698] = 32'he44a929e;
    ram_cell[     699] = 32'h7c439f8e;
    ram_cell[     700] = 32'hed808a53;
    ram_cell[     701] = 32'h62b3005f;
    ram_cell[     702] = 32'hd3c22cda;
    ram_cell[     703] = 32'h50cb2755;
    ram_cell[     704] = 32'h1c64c0ca;
    ram_cell[     705] = 32'h65779b74;
    ram_cell[     706] = 32'hb6cc3285;
    ram_cell[     707] = 32'ha3028386;
    ram_cell[     708] = 32'h117a7d4f;
    ram_cell[     709] = 32'ha5858b7b;
    ram_cell[     710] = 32'h31ebcc43;
    ram_cell[     711] = 32'h4fa52726;
    ram_cell[     712] = 32'hcd6025e2;
    ram_cell[     713] = 32'ha33d5290;
    ram_cell[     714] = 32'h382a0250;
    ram_cell[     715] = 32'h6a5c5925;
    ram_cell[     716] = 32'h6d50a3be;
    ram_cell[     717] = 32'hbb6a1a29;
    ram_cell[     718] = 32'hcdb251c4;
    ram_cell[     719] = 32'hd5a33248;
    ram_cell[     720] = 32'hc484e3e2;
    ram_cell[     721] = 32'h7a2a1cf8;
    ram_cell[     722] = 32'h9b2d42ec;
    ram_cell[     723] = 32'h0caddf6b;
    ram_cell[     724] = 32'h1982ee82;
    ram_cell[     725] = 32'h9eb0de06;
    ram_cell[     726] = 32'h17295ad9;
    ram_cell[     727] = 32'ha7c8d305;
    ram_cell[     728] = 32'ha1b8ecc8;
    ram_cell[     729] = 32'h1d8664a8;
    ram_cell[     730] = 32'h5343c376;
    ram_cell[     731] = 32'hf5c87a04;
    ram_cell[     732] = 32'hedde9cea;
    ram_cell[     733] = 32'hcadc07e7;
    ram_cell[     734] = 32'hf44e51af;
    ram_cell[     735] = 32'hf38556e7;
    ram_cell[     736] = 32'hc140f734;
    ram_cell[     737] = 32'h11fc0a15;
    ram_cell[     738] = 32'h11b21917;
    ram_cell[     739] = 32'h91cebb27;
    ram_cell[     740] = 32'h22344f12;
    ram_cell[     741] = 32'h161cd5dc;
    ram_cell[     742] = 32'hb5e95137;
    ram_cell[     743] = 32'h3e3c4bdb;
    ram_cell[     744] = 32'h8414c0b6;
    ram_cell[     745] = 32'hd160c990;
    ram_cell[     746] = 32'hea887baa;
    ram_cell[     747] = 32'h048f6319;
    ram_cell[     748] = 32'hb17cdc09;
    ram_cell[     749] = 32'h17ef4306;
    ram_cell[     750] = 32'h92fef17b;
    ram_cell[     751] = 32'h219d8a81;
    ram_cell[     752] = 32'hffad0d12;
    ram_cell[     753] = 32'h5ee5c7d4;
    ram_cell[     754] = 32'hbf9186a9;
    ram_cell[     755] = 32'hd6b6369e;
    ram_cell[     756] = 32'hcb2d4e9f;
    ram_cell[     757] = 32'h4fb3757b;
    ram_cell[     758] = 32'h395d2676;
    ram_cell[     759] = 32'h16d50318;
    ram_cell[     760] = 32'h6e16b572;
    ram_cell[     761] = 32'h17e2a566;
    ram_cell[     762] = 32'hd2c4af2d;
    ram_cell[     763] = 32'h10a13b42;
    ram_cell[     764] = 32'h404a0c92;
    ram_cell[     765] = 32'hfc0a0642;
    ram_cell[     766] = 32'h15c6bfdf;
    ram_cell[     767] = 32'hc17f7ed5;
end

endmodule

